Inverter Simulation

* this file edited to remove everything not ion tt lib
.lib "/home/sandman/pdks/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* instantiate inverter
Xinv Y A VPWR VGND VPWR inverter

.subckt inverter Y A NWELL VSUBS VGND VPWR
X0 Y A VPWR NWELL sky130_fd_pr__pfet_01v8 ad=5.5e+11p pd=3.1e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 Y A VGND SUB sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=2.4e+06u as=2.3e+11p ps=2.3e+06u w=650000u l=150000u
.ends

* set GND and PWR
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00

.control
run
plot A Y
.endc

.end
